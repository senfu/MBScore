`resetall
module MBScore_rf(
    
);